    Mac OS X            	   2   �      �                                      ATTR       �   �   =                  �     com.apple.TextEncoding      �   .  com.dropbox.attributes   utf-8;134217984x��V*�/άP�R�VJ�HM.-IL�IsSK�%�@[[���Z @